library ieee;
use ieee.std_logic_1164.all;
use work.arch_defs.all;

entity memoryAccess is
    port();
end;

architecture struct of memoryAccess is



begin



end struct;
