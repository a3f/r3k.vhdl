library ieee;
use ieee.std_logic_1164.all;
use work.arch_defs.all;

entity memoryAccess is
    port(
	ALUResult, regReadData2 : in word_t;
	signExtend : in ctrl_t);
end;

architecture struct of memoryAccess is



begin

	

end struct;
