-- SKIP Tests regfile, ALU and related MUXes/Extenders
